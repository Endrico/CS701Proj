library ieee;
use ieee.std_logic_1164.all; 

ENTITY register_32 is port(
	clk	:	in	std_logic;
	enable:	in	std_logic;
	reset	:	in std_logic;
	input	:	in std_logic_vector(31 downto 0);
	output:	out std_logic_vector(31 downto 0)
	
);
END register_32;

architecture behaviour of register_32 is
begin 
	process(clk)
		begin
			if (clk = '1' and clk'event) then
				if (reset = '1') then
					output <= x"00000000";  -- x stands for hexidecimal 16 bits long  therefor four zeros
				elsif (enable = '1') then
					output <= input;
				end if;
			end if;
	end process;
end behaviour; 

