library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
use IEEE.NUMERIC_STD.ALL;

ENTITY MAX IS
	PORT
	(
		A, B : IN STD_LOGIC_VECTOR(15 downto 0);
		max_out : OUT STD_LOGIC_VECTOR(15 downto 0)
	);
END MAX;

ARCHITECTURE bhvr OF MAX IS
BEGIN
	max_out <= A when A > B else
			   B;
end ARCHITECTURE bhvr;

