library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity test_bench is 
end test_bench;

architecture behaviour of test_bench is 
	component processor
	
	port(
			-- place the stuff for the processor here all processor ports	
			
		 );
	end component;
	